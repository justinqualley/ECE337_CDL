// $Id: $
// File name:   encoder.sv
// Created:     4/27/2022
// Author:      Robert Sego
// Lab Section: 337-015
// Version:     1.0  Initial Design Entry
// Description: encoder

module encoder (



);

endmodule